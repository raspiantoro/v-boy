module config

pub const(
	pixel_width = 160
	pixel_height = 144
)